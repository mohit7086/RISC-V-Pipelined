module name(
    input clk,
    input rst,
    input [31:0] PC,
    

);
    
endmodule